LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY adder_tree IS
	GENERIC (

	);
	PORT (

	);
END adder_tree;

ARCHITECTURE Behavioral OF adder_tree IS

BEGIN

END Behavioral;